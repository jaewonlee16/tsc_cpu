module cache
   (
    input clk,
    input reset_n,
    input read_cache,
    input write_cache,
    input [WORD_SIZE-1:0] address_cache,
    inout [WORD_SIZE-1:0] data_cache_datapath, // data connected to datapath
    inout [4 * READ_SIZE - 1 : 0] data_mem_cache, // data connected to memory

    output doneWrite,  // tells the cpu that writing is finshed
    output [WORD_SIZE-1:0] address_memory,
    output readM,
    output writeM,
   );
    reg [`WORD_SIZE-1:0] temp_data;
    reg [`WORD_SIZE-1:0] num_cache_access,    // for debugging
    reg [`WORD_SIZE-1:0] num_cache_miss,      // for debugging

   // for data_cache_datapath
    reg [`WORD_SIZE - 1 : 0] cache_output_data;
    reg [4 * `WORD_SIZE - 1 : 0] mem_output_data;


    // 4 line, 4 word wide cache block
    // as line number is 4, index is log(4) = 2 bits
    // as block size is 4, block offset is log(4) = 2bits
    // therefore, tag is 16 - 2 - 2 = 12 bits
    reg [4*`WORD_SIZE-1:0]  data_bank[3:0];
    reg [`WORD_SIZE-5:0]    tag_bank[3:0];
    reg [3:0]              valid;

   // Address decoding
   wire [1:0] index;
   wire [`WORD_SIZE-5:0] tag;
   wire [1:0] block_offset;             
   assign index = address_cache[3:2];
   assign tag = address_cache[`WORD_SIZE-1:4];
   assign block_offset = address_cache[1:0];

   // data_bank decoding
   wire [`WORD_SIZE - 1:0] block_0;  // block offset 0
   wire [`WORD_SIZE - 1:0] block_1;  // block offset 1
   wire [`WORD_SIZE - 1:0] block_2;  // block offset 2
   wire [`WORD_SIZE - 1:0] block_3;  // block offset 3
   
   assign {block_0, block_1, block_2, block_3} = data_bank[index];

   // ouput port assignment
   assign data_mem_cache = writeM ? mem_output_data : 4*`WORD_SIZE'bz;
   assign data_cache_datapath = read_cache ? cache_output_data : `WORD_SIZE'bz;


   // cache hit
   wire hit;
   assign hit = valid[index] && (tag_bank[index] == tag) 
               && data_bank[index] [63 : 60] != `OPCODE_NOP;

   // memory signals
   assign readM = (read_cache || write_cache) && !hit;


   always @ (*) begin
      if (read_cache && !hit) begin

      end
   end

   always @ (posedge clk) begin
      if (!reset_n) begin
         for (i=0; i<4; i=i+1) begin
            data_bank[i] <= 0;
            tag_bank[i] <= 0;
            valid[i] <= 0;
            dirty[i] <= 0;
            num_cache_miss <= 0;
            num_cache_access <= 0;

         end
      end
      else begin
         // Request type: Read
         if (read_cache) begin
            if (!hit) begin
               // Read data from lower memory into the cache block
               data_bank[index] <= data_mem_cache;
               readM <= 1;
            end
            else readM <= 0;
             

         end
         // Request type : Write
         else if (write_cache) begin
            if (!hit) begin
               // Read data from lower memory into the cache block
               data_bank[index] <= data_mem_cache;
               readM <= 1;
            end
            else readM <= 0;

         end
         // Request type: No memory request
         else begin

         end 
      end
   end